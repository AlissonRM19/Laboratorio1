module Processor ();

endmodule